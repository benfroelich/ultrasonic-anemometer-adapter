* HCMOS Subcircuit and Primitive Elements Library
* hc_tfast.cir
* Fast Process Corner
* Standard Logic Product Group
* NXP Semiconductors
*
* Version Date       By   Remarks
* ---------------------------------------------------------------------
*    1.2  30/03/2011 RRV  Rewritten netlists to add package options.
*    1.12 27/10/2010 RRV  Added HC(T)240/253
*    1.11 06/07/2010 RRV  Added HC(T)02/08/86
*    1.10 10/12/2009 RRV  Removed HCT05
*    1.09 09/22/2009 RRV  Corrected typo in SWITCH3N
*    1.08 09/08/2009 RRV  Added HC(T)4020/4060
*    1.07 03/27/2009 RRV  Added HC(T)05
*    1.06 02/20/2006 RRV  Added HC(T)366/368
*    1.05 10/27/2005 RRV  Updated HC/T04 and HCU04 models
*    1.04 09/22/2003 RM   Active High Enable for SWI2 and SWI2T
*
************************************************
*           FAST N-Channel Transistor          *
*            UCB-3 Parameter Set               *
*         HIGH-SPEED CMOS Logic Family         *
*                10-Jan.-1995                  *
************************************************
.Model MHCNEF NMOS
+LEVEL = 3
+KP    = 49.6E-6
+VTO   = 0.52
+TOX   = 49.0E-9
+NSUB  = 4.0E15
+GAMMA = 0.74
+PHI   = 0.65
+VMAX  = 135E3
+RS    = 30
+RD    = 30
+XJ    = 0.10E-6
+LD    = 0.69E-6
+DELTA = 0.38
+THETA = 0.048
+ETA   = 0.020
+KAPPA = 0.0
+WD    = 0.5E-6

***********************************************
*          FAST P-Channel transistor          *
*           UCB-3 Parameter Set               *
*         HIGH-SPEED CMOS Logic Family        *
*                10-Jan.-1995                 *
***********************************************
.Model MHCPEF PMOS
+LEVEL = 3
+KP    = 24.6E-6
+VTO   = -0.51
+TOX   = 49.0E-9
+NSUB  = 3.6E16
+GAMMA = 0.82
+PHI   = 0.65
+VMAX  = 600E3
+RS    = 60
+RD    = 60
+XJ    = 0.61E-6
+LD    = 0.35E-6
+DELTA = 2.12
+THETA = 0.100
+ETA   = 0.260
+KAPPA = 0.0
+WD    = 0.5E-6


.MODEL  INT D


****************************************
*   START OF SUB-CIRCUIT DESCRIPTION   *
*            MARCH 30, 2011            *
****************************************

*****NOMIN.CIR*****

****Version 1.04 Added Inverter****
.SUBCKT INV4F    2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
MP1 3  2 50 50  MHCPEF W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2 60 60  MHCNEF W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
.ENDS


.SUBCKT INP0F   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  3  100
MP1 3 50 50 50  MHCPEF W=20U L=2.4U AD=100P AS=100P PD=40U PS= 20U
MN1 3 60 60 60  MHCNEF W=35U L=2.4U AD=260P AS=260P PD=70U PS= 20U
.ENDS

.SUBCKT INP1F   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEF W=20U L=2.4U AD=100P AS=100P PD=40U PS= 20U
MN1 4 60 60 60  MHCNEF W=35U L=2.4U AD=260P AS=260P PD=70U PS= 20U
MP2 3  4 50 50  MHCPEF W=88U L=2.4U AD=290P AS=550P PD=10U PS=100U
MN2 3  4 60 60  MHCNEF W=56U L=2.4U AD=162P AS=550P PD=10U PS= 75U
.ENDS

.SUBCKT INP1TF   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEF W= 20U L=2.4U AD=100P AS=100P PD= 40U PS= 20U
MN1 4 60 60 60  MHCNEF W= 35U L=2.4U AD=260P AS=260P PD= 70U PS= 20U
MP2 3  4  5 50  MHCPEF W= 88U L=2.4U AD=290P AS=550P PD=107U PS=195U
MN2 3  4 60 60  MHCNEF W= 56U L=2.4U AD=162P AS=550P PD= 55U PS=162U
D1 50  5  INT
MP4 3  6 50 50  MHCPEF W=6.4U L=4.0U AD= 60P AS= 60P PD=13U PS= 24U
MN4 3  4 60 60  MHCNEF W=185U L=2.4U AD=740P AS=740P PD=50U PS=185U
MP5 6  3 50 50  MHCPEF W=6.4U L=3.2U AD= 50P AS= 50P PD=10U PS= 20U
MN5 6  3 60 60  MHCNEF W=6.4U L=3.2U AD= 50P AS= 50P PD=10U PS= 20U
.ENDS

.SUBCKT INP2F   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEF W= 20U L=2.4U AD=100P AS=100P PD=40U PS= 20U
MN1 4 60 60 60  MHCNEF W= 35U L=2.4U AD=260P AS=260P PD=70U PS= 20U
MP2 3  4 50 50  MHCPEF W=176U L=2.4U AD=580P AS=580P PD=10U PS=200U
MN2 3  4 60 60  MHCNEF W=112U L=2.4U AD=325P AS=580P PD=10U PS=150U
.ENDS

.SUBCKT INP2TF   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEF W= 20U L=2.4U AD=100P AS= 100P PD=40U PS= 20U
MN1 4 60 60 60  MHCNEF W= 35U L=2.4U AD=260P AS= 260P PD=70U PS= 20U
MP2 3  4  5 50  MHCPEF W=176U L=2.4U AD=580P AS=1100P PD=10U PS=200U
MN2 3  4 60 60  MHCNEF W=112U L=2.4U AD=325P AS=1100P PD=10U PS=150U
D1 50  5   INT
MP4 3  6 50 50  MHCPEF W=6.4U L=4.0U AD= 60P AS= 60P PD=13U PS= 24U
MN4 3  4 60 60  MHCNEF W=348U L=2.4U AD=740P AS=740P PD=50U PS=348U
MP5 6  3 50 50  MHCPEF W=6.4U L=3.2U AD= 50P AS= 50P PD=10U PS= 20U
MN5 6  3 60 60  MHCNEF W=6.4U L=3.2U AD= 50P AS= 50P PD=10U PS= 20U
.ENDS


.SUBCKT SMT1F   2  3  50  60
* SCHMITT-TRIGGER INPUT FOR HC14 CMOS INPUT LEVELS
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEF W=20U L=2.4U AD=100P AS=100P PD=40U PS=20U
MN1 4 60 60 60  MHCNEF W=35U L=2.4U AD=140P AS=140P PD=50U PS=35U
MP2 5  4 50 50  MHCPEF W=36U L=2.4U AD=140P AS=140P PD=50U PS=35U
MN2 6  4 60 60  MHCNEF W=16U L=2.4U AD= 70P AS= 70P PD=15U PS=17U
MP3 3  4  5 50  MHCPEF W=44U L=2.4U AD=220P AS=220P PD=60U PS=44U
MN3 3  4  6  6  MHCNEF W=17U L=2.4U AD= 70P AS= 70P PD=15U PS=16U
MP4 5  3 60 50  MHCPEF W=36U L=2.4U AD=150P AS=150P PD=60U PS=36U
MN4 6  3 50  6  MHCNEF W= 6U L=  4U AD= 25P AS= 25P PD=10U PS= 6U
.ENDS


.SUBCKT SMTTL1F   2  3  50  60
* SCHMITT-TRIGGER INPUT FOR HCT14 WITH TTL INPUT LEVELS
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEF W= 20U L=2.4U AD= 100P AS= 100P PD= 40U PS= 20U
MN1 4 60 60 60  MHCNEF W= 35U L=2.4U AD= 140P AS= 140P PD= 50U PS= 35U
D1  50  7  INT
MP2 5  4  7  7  MHCPEF W= 36U L=2.4U AD= 140P AS= 140P PD= 50U PS= 35U
MN2 6  4 60 60  MHCNEF W=216U L=2.4U AD= 860P AS= 860P PD=140U PS=216U
MP3 3  4  5 50  MHCPEF W= 54U L=2.4U AD= 220P AS= 220P PD= 60U PS= 44U
MN3 3  4  6  6  MHCNEF W=257U L=2.4U AD=1000P AS=1000P PD=150U PS=257U
MP4 5  3 60 50  MHCPEF W= 32U L=  4U AD= 120P AS= 120P PD=100U PS= 32U
MN4 6  3 50  6  MHCNEF W= 14U L=  4U AD= 100P AS= 100P PD= 30U PS= 24U
MP5 8  3 50 50  MHCPEF W= 10U L=2.4U AD=  40P AS=  40P PD= 16U PS= 10U
MN5 8  3 60 60  MHCNEF W=  5U L=2.4U AD=  20P AS=  20P PD= 12U PS=  5U
MP6 3  8 50 50  MHCPEF W=  6U L=8.0U AD=  30P AS=  30P PD= 16U PS=  6U
.ENDS


.SUBCKT INVF    2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
MP1 3  2 50 50  MHCPEF W=364U L=2.4U AD=500P  AS=500P PD=10U PS=430U
MN1 3  2 60 60  MHCNEF W=184U L=2.4U AD=275P  AS=275P PD=10U PS=270U
.ENDS


.SUBCKT NANDF   2  3  4  50  60
*INTERNAL NAND
*IN1 = 2, IN2 = 3, OUT = 4, VCC= 50, GND = 60
MP1 4  2  50  50  MHCPEF W=112U  L=2.4U AD=150P AS=300P PD= 75U PS=150U
MP2 4  3  50  50  MHCPEF W=112U  L=2.4U AD=150P AS=300P PD= 75U PS=150U
MN1 4  2   5  60  MHCNEF W=300U  L=2.4U AD=300P AS=300P PD=300U PS=300U
MN2 5  3  60  60  MHCNEF W=300U  L=2.4U AD=300P AS=300P PD=300U PS=300U
.ENDS


.SUBCKT LLCF   2  3  40  50  60
* LEVEL CONVERTER
* INA = 2,  OUT = 3,  VEE = 40,  VCC = 50,  GND =  60
MP4 4  2  50  50  MHCPEF W= 30U  L= 2.4U AD=120P AS=120P PD= 40U PS= 30U
MN4 4  2  60  60  MHCNEF W= 15U  L= 2.4U AD= 60P AS= 60P PD= 20U PS= 15U
MP1 5  4  50  50  MHCPEF W=135U  L= 2.4U AD=500P AS=500P PD=100U PS=135U
MP2 6  2  50  50  MHCPEF W=135U  L= 2.4U AD=500P AS=500P PD=100U PS=135U
MN1 5  6  40  40  MHCNEF W=6.4U  L=18.8U AD= 25P AS= 25P PD= 20U PS=6.4U
MN2 6  5  40  40  MHCNEF W=6.4U  L=18.8U AD= 25P AS= 25P PD= 20U PS=6.4U
MP3 7  6  50  50  MHCPEF W= 10U  L= 4.0U AD= 40P AS= 40P PD= 20U PS= 10U
MN3 7  6  40  40  MHCNEF W=  5U  L= 4.0U AD= 20P AS= 20P PD= 10U PS=  5U
MP5 3  7  50  50  MHCPEF W= 30U  L= 2.4U AD=120P AS=120P PD= 40U PS= 30U
MN5 3  7  40  40  MHCNEF W= 15U  L= 2.4U AD= 60P AS= 60P PD= 20U PS= 15U
.ENDS

.SUBCKT SWITCH1F   2  8  9  40  50
* ANALOG SWITCH
* INPUT = 2,   Y = 8,  Z = 9,  VEE = 40,  VCC =50
MP1 3  2  50  50  MHCPEF W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2  40  40  MHCNEF W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
MP4 4  3  50  50  MHCPEF W= 350U L=2.4U AD= 900P AS= 900P PD=200U PS= 350U
MN4 4  3  40  40  MHCNEF W= 150U L=2.4U AD= 400P AS= 400P PD=100U PS= 150U
MP5 8  4   5  50  MHCPEF W= 216U L=2.4U AD= 900P AS= 900P PD=100U PS= 216U
MN5 8  3   5   5  MHCNEF W= 108U L=2.4U AD= 430P AS= 430P PD= 50U PS= 108U
MN6 5  4  40  40  MHCNEF W= 145U L=2.4U AD= 600P AS= 600P PD= 75U PS= 145U
MP7 9  4   8  50  MHCPEF W=1068U L=2.4U AD=2500P AS=2500P PD= 10U PS=1068U
MN7 9  3   8   5  MHCNEF W= 312U L=2.4U AD=1200P AS=1200P PD= 10U PS= 312U
.ENDS

.SUBCKT SWITCH2F   2  8  9  50  60
* ANALOG SWITCH
* INPUT= 2   Y= 8   Z= 9  VCC= 50   GND= 60
MP1 3  2  50  50  MHCPEF W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2  60  60  MHCNEF W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
MP4 4  3  50  50  MHCPEF W= 350U L=2.4U AD= 900P AS= 900P PD=200U PS= 350U
MN4 4  3  60  60  MHCNEF W= 150U L=2.4U AD= 400P AS= 400P PD=100U PS= 150U
MP5 5  3   8  50  MHCPEF W=  85U L=2.4U AD= 355P AS= 355P PD= 40U PS=  85U
MN5 5  4   8   5  MHCNEF W=  42U L=2.4U AD= 170P AS= 170P PD= 20U PS=  42U
MN6 5  3  60  60  MHCNEF W= 145U L=2.4U AD= 600P AS= 600P PD= 75U PS= 145U
MP7 9  3   8  50  MHCPEF W=1900U L=2.4U AD=2500P AS=2500P PD= 10U PS=1900U
MN7 9  4   8   5  MHCNEF W= 576U L=2.4U AD=1200P AS=1200P PD= 10U PS= 576U
.ENDS

.SUBCKT SWITCH3F   2  8  9  40  50
* ANALOG SWITCH
* INPUT = 2   Y = 8  Z = 9  VEE = 40  VCC = 50
MP1 3  2  50  50  MHCPEF W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2  40  40  MHCNEF W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
MP4 4  3  50  50  MHCPEF W= 350U L=2.4U AD= 900P AS= 900P PD=200U PS= 350U
MN4 4  3  40  40  MHCNEF W= 150U L=2.4U AD= 400P AS= 400P PD=100U PS= 150U
MP5 9  3   8  50  MHCPEF W=1168U L=2.4U AD=2730P AS=2730P PD= 10U PS=1168U
MN5 9  4   8  40  MHCNEF W= 312U L=2.4U AD=1200P AS=1200P PD= 10U PS= 312U
.ENDS


.SUBCKT BUSOUTPF   2   3   4   50   60
* INPUT = 2  OEN = 3 (LOW)  OUT = 4  VCC = 50  GND = 60
* 3-STATE BUS OUTPUT
MP1 5  3   50  50  MHCPEF W= 90U  L=2.4U AD= 360P AS= 360P PD= 30U PS=360U
MN1 5  3   60  60  MHCNEF W= 40U  L=2.4U AD= 160P AS= 160P PD= 20U PS= 40U
MP2 6  2   50  50  MHCPEF W=480U  L=2.4U AD=1800P AS=1800P PD=100U PS=480U
MN2 7  2   60  60  MHCNEF W=240U  L=2.4U AD=1000P AS=1000P PD= 50U PS=240U
MP3 7  3    6  50  MHCPEF W=280U  L=2.4U AD=1120P AS=1120P PD= 55U PS=280U
MN3 7  3   60  60  MHCNEF W=160U  L=2.4U AD= 640P AS= 640P PD= 40U PS=160U
MP4 6  5   50  50  MHCPEF W=240U  L=2.4U AD=1000P AS=1000P PD= 50U PS=240U
MN4 7  5    7  60  MHCNEF W=190U  L=2.4U AD= 760P AS= 760P PD= 45U PS=190U
R1  6  8  200
R2  7  9  200
MP5 4  8   50  50  MHCPEF W=540U  L=2.4U AD=1500P AS=1500P PD=10U PS=540U
MN5 4  9   60  60  MHCNEF W=233U  L=2.4U AD= 750P AS= 750P PD=10U PS=233U
R3  8  10 100
R4  9  11 100
MP6 4  10  50  50  MHCPEF W=540U  L=2.4U AD=1500P AS=1500P PD=10U PS=540U
MN6 4  11  60  60  MHCNEF W=233U  L=2.4U AD= 750P AS= 750P PD=10U PS=233U
R5 10  12  50
R6 11  13  50
MP7 4  12  50  50  MHCPEF W=540U  L=2.4U AD=1500P AS=1500P PD=10U PS=540U
MN7 4  13  60  60  MHCNEF W=233U  L=2.4U AD= 750P AS= 750P PD=10U PS=233U
.ENDS

.SUBCKT OUTUF  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2 4 100
MP1 3 4 50 50  MHCPEF W=485U L=2.4U AD=1200P AS=530P PD=10U PS=180U
MN1 3 4 60 60  MHCNEF W=222U L=2.4U AD=530P AS=300P PD=10U PS=130U
R2  4 5 50
MP2 3 5 50 50  MHCPEF W=485U L=2.4U AD=1200P AS=530P PD=10U PS=180U
MN2 3 5 60 60  MHCNEF W=222U L=2.4U AD=530P AS=300P PD=10U PS=130U
R3  5 6 50
MP3 3 6 50 50  MHCPEF W=485U L=2.4U AD=1200P AS=530P PD=10U PS=180U
MN3 3 6 60 60  MHCNEF W=222U L=2.4U AD=530P AS=300P PD=10U PS=130U
.ENDS

.SUBCKT OUTPF  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2 4 100
MP1 3 4 50 50  MHCPEF W=360U L=2.4U AD=400P AS=400P PD=10U PS=180U
MN1 3 4 60 60  MHCNEF W=140U L=2.4U AD=200P AS=300P PD=10U PS=130U
R2  4 5 50
MP2 3 5 50 50  MHCPEF W=360U L=2.4U AD=400P AS=400P PD=10U PS=180U
MN2 3 5 60 60  MHCNEF W=140U L=2.4U AD=200P AS=200P PD=10U PS=130U
R3  5 6 50
MP3 3 6 50 50  MHCPEF W=360U L=2.4U AD=400P AS=400P PD=10U PS=180U
MN3 3 6 60 60  MHCNEF W=140U L=2.4U AD=200P AS=200P PD=10U PS=130U
.ENDS

.SUBCKT OUTPODF  2  3  60
*IN=2, OUT=3, GND=60
R1  2 4 50
MN1 3 4 60 60  MHCNEF W=140U L=2.4U AD=200P AS=300P PD=10U PS=130U
R2  4 5 25
MN2 3 5 60 60  MHCNEF W=140U L=2.4U AD=200P AS=200P PD=10U PS=130U
R3  5 6 25
MN3 3 6 60 60  MHCNEF W=140U L=2.4U AD=200P AS=200P PD=10U PS=130U
.ENDS

.SUBCKT INPOSCF   2  5  3  50  60
R1  2  4  100
MP1 4 50 50 50  MHCPEF W=20U  L=2.4U AD=100P AS=100P PD=40U PS=20U
MN1 4 60 60 60  MHCNEF W=35U  L=2.4U AD=260P AS=260P PD=70U PS=20U
MP2 6  4 50 50  MHCPEF W=707U L=2.4U AD=1700P AS=2000P PD=40U PS=60U
MP3 6  5 50 50  MHCPEF W=166U L=2.4U AD=400P AS=800P PD=40U PS=60U
MN2 6  4  7 60  MHCNEF W=480U L=2.4U AD=1200P AS=900P PD=60U PS=65U
MN3 7  5 60 60  MHCNEF W=640U L=2.4U AD=1200P AS=2000P PD=90U PS=80U
MP4 3  6 50 50  MHCPEF W=832U L=2.4U AD=2000P AS=3000P PD=40U PS=60U
MN4 3  6 60 60  MHCNEF W=333U L=2.4U AD=800P AS=1600P PD=40U PS=60U
.ENDS

.SUBCKT INP3F   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEF W=20U  L=2.4U AD=100P AS=100P PD=40U PS=20U
MN1 4 60 60 60  MHCNEF W=35U  L=2.4U AD=260P AS=260P PD=70U PS=20U
MP2 5  4 50 50  MHCPEF W=29U  L=2.4U AD=85P AS=85P PD=29U PS=29U
MN2 5  4 60 60  MHCNEF W=19U  L=2.4U AD=70P AS=70P PD=19U PS=19U
MP3 3  5 50 50  MHCPEF W=112U L=2.4U AD=200P AS=200P PD=30U PS=30U
MN3 3  5 60 60  MHCNEF W=56U  L=2.4U AD=100P AS=100P PD=15U PS=15U
.ENDS

.SUBCKT INP3TF   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEF W=20U  L=2.4U AD=100P AS=100P PD=40U PS=20U
MN1 4 60 60 60  MHCNEF W=35U  L=2.4U AD=260P AS=260P PD=70U PS=20U
MP2 6  4  5 50  MHCPEF W=29U  L=2.4U AD=85P AS=85P PD=29U PS=29U
MN2 6  4 60 60  MHCNEF W=19U  L=2.4U AD=70P AS=70P PD=19U PS=19U
D1 50  5   INT
MP4 6  3 50 50  MHCPEF W=6.4U L=4.0U AD=25P AS=25P PD=6.4U PS=6.4U
MN4 6  4 60 60  MHCNEF W=80U  L=2.4U AD=120P AS=240P PD=80U PS=80U
MP5 3  6 50 50  MHCPEF W=112U L=3.2U AD=200P AS=200P PD=30U PS=30U
MN5 3  6 60 60  MHCNEF W=56U  L=3.2U AD=100P AS=100P PD=15U PS=15U
.ENDS
*******************************************************************
*******************************************************************

******CIR_NOMIN-HC TYPES******

.SUBCKT INV0  20 30 80 90
*IN=20, OUT=30, VCC=80, GND=90
XINP  20  25  80  90    INP0F
XOUTP 25  30  80  90    OUTUF
.ENDS


.SUBCKT INV1  20 30 80 90
*IN=20, OUT=30, VCC=80, GND=90
XINP  20  25  80  90    INP1F
XINV  25  35  80  90    INVF
XOUTP 35  30  80  90    OUTPF
.ENDS


.SUBCKT INV2  20  30  80 90
*IN=20, OUT=30, VCC=80, GND=90
XINP  20  25  80  90    INP2F
XINV  25  35  80  90    INVF
XOUTP 35  30  80  90    OUTPF
.ENDS

.SUBCKT INVOD  20  30  80  90
*IN=20, OUT=30, VCC=80, GND=90
XINP    20  25  80  90    INP2F
XINV    25  35  80  90    INVF
XOUTPOD 35  30  90        OUTPODF
.ENDS

.SUBCKT INVSMT  20  30  80 90
*IN=20, OUT=30, VCC=80, GND=90
XINP  20  25  80  90    SMT1F
XINV  25  35  80  90    INVF
XOUTP 35  30  80  90    OUTPF
.ENDS

.SUBCKT NINV1  20  30  80 90
*IN=20, OUT=30, VCC=80, GND=90
XINP  20  25  80  90    INP1F
XINV0 25  35  80  90    INVF
XINV1 35  45  80  90    INVF
XOUTP 45  30  80  90    OUTPF
.ENDS

.SUBCKT NANDINV 20  50  30  80  90
*INVERTING 2-NAND
*EN = 50, IN = 20, OUT = 30, VCC = 80, GND = 90
XIN1  20  25      80  90   INP2F
XIN2  50  35      80  90   INP2F
XNAND 25  35  36  80  90   NANDF
XOUT  36  30      80  90   OUTPF
.ENDS

.SUBCKT SWI1  20  30  40  70  80  90
* INP = 20  Y = 30  Z = 40  VEE = 70  VCC = 80  GND = 90
XINP 20  25  80  90      INP2F
XLC  25  35  70  80  90  LLCF
XAS  35  30  40  70  80  SWITCH1F
.ENDS


.SUBCKT SWI2  20 30 40 80 90
* INP = 20 Y = 30 Z = 40 VCC = 80  GND = 90
*XINP  20  25  80  90      INP2F
****Version 1.04 Inserted inverter****
XINP  20  250      80  90  INP2F
XINV  250  25      80  90  INV4F
XAS   25   30  40  80  90  SWITCH2F
.ENDS


.SUBCKT SWI3  20  30  40  70  80  90
* INP = 20  Y = 30  Z = 40  VEE = 70  VCC = 80  GND = 90
XINP 20  25  80  90      INP1F
XLC  25  35  70  80  90  LLCF
XAS  35  30  40  70  80  SWITCH3F
.ENDS


.SUBCKT NINV3  20  50  30  80  90
* INP = 20  OEN = 50(LOW)  OUT = 30   VCC = 80  GND = 90
XINP      20  25  80  90      INP2F
XINV      25  35  80  90      INVF
XBUSOUTP  35  50  30  80  90  BUSOUTPF
.ENDS

.SUBCKT INV3  20  50  30  80  90
* INP = 20  OEN = 50(LOW)  OUT = 30   VCC = 80  GND = 90
XINP      20  25  80  90      INP2F
XBUSOUTP  25  50  30  80  90  BUSOUTPF
.ENDS

.SUBCKT OSC  20  50  30  80  90
*
* INP = 20  MR = 50  OUT = 30  VCC = 80  GND = 90
XINPOSC   20  17  25  80  90  INPOSCF
XINV1     25  35  80  90      INVF
XOUTPN    35  30  80  90      OUTPF
XINPMR	  50  16  80  90      INP3F
XINV2     16  17  80  90      INVF
.ENDS

******CIR_NOMIN-HCT TYPES******

.SUBCKT INV1T  20 30 80 90
*IN=20, OUT=30, VCC=80, GND=90
XINP  20  25  80  90    INP1TF
XINV  25  35  80  90    INVF
XOUTP 35  30  80  90    OUTPF
.ENDS


.SUBCKT INV2T  20  30  80 90
*IN=20, OUT=30, VCC=80, GND=90
XINP  20  25  80  90    INP2TF
XINV  25  35  80  90    INVF
XOUTP 35  30  80  90    OUTPF
.ENDS

.SUBCKT INVODT  20  30  80  90
*IN=20, OUT=30, VCC=80, GND=90
XINP    20  25  80  90    INP2TF
XINV    25  35  80  90    INVF
XOUTPOD 35  30  90        OUTPODF
.ENDS

.SUBCKT INVSMTT  20  30  80 90
*IN=20, OUT=30, VCC=80, GND=90
XINP  20  25  80  90    SMTTL1F
XINV  25  35  80  90    INVF
XOUTP 35  30  80  90    OUTPF
.ENDS

.SUBCKT NINV1T  20  30  80 90
*IN=20, OUT=30, VCC=80, GND=90
XINP  20  25  80  90    INP1TF
XINV0 25  35  80  90    INVF
XINV1 35  45  80  90    INVF
XOUTP 45  30  80  90    OUTPF
.ENDS

.SUBCKT NANDINVT 20  50  30  80  90
*INVERTING 2-NAND
*EN = 50, IN = 20, OUT = 30, VCC = 80, GND = 90
XIN1  20  25      80  90   INP2TF
XIN2  50  35      80  90   INP2TF
XNAND 25  35  36  80  90   NANDF
XOUT  36  30      80  90   OUTPF
.ENDS

.SUBCKT SWI1T  20  30  40  70  80  90
* INP = 20  Y = 30  Z = 40  VEE = 70  VCC = 80  GND = 90
XINP 20  25  80  90      INP2TF
XLC  25  35  70  80  90  LLCF
XAS  35  30  40  70  80  SWITCH1F
.ENDS


.SUBCKT SWI2T  20 30 40 80 90
* INP = 20 Y = 30 Z = 40 VCC = 80  GND = 90
*XINP  20  25  80  90      INP2TF
****Version 1.04 Inserted inverter****
XINP  20  250      80  90  INP2TF
XINV  250  25      80  90  INV4F
XAS   25   30  40  80  90  SWITCH2F
.ENDS


.SUBCKT SWI3T  20  30  40  70  80  90
* INP = 20  Y = 30  Z = 40  VEE = 70  VCC = 80  GND = 90
XINP 20  25  80  90      INP1TF
XLC  25  35  70  80  90  LLCF
XAS  35  30  40  70  80  SWITCH3F
.ENDS


.SUBCKT NINV3T  20  50  30  80  90
* INP = 20  OEN = 50(LOW)  OUT = 30   VCC = 80  GND = 90
XINP      20  25  80  90      INP2TF
XINV      25  35  80  90      INVF
XBUSOUTP  35  50  30  80  90  BUSOUTPF
.ENDS

.SUBCKT INV3T  20  50  30  80  90
* INP = 20  OEN = 50(LOW)  OUT = 30   VCC = 80  GND = 90
XINP      20  25  80  90      INP2TF
XBUSOUTP  25  50  30  80  90  BUSOUTPF
.ENDS

.SUBCKT OSCT  20  50  30  80  90
*
* INP = 20  MR = 50  OUT = 30  VCC = 80  GND = 90
XINPOSC   20  17  25  80  90  INPOSCF
XINV1     25  35  80  90      INVF
XOUTPN    35  30  80  90      OUTPF
XINPMR	  50  16  80  90      INP3TF
XINV2     16  17  80  90      INVF
.ENDS

***********************************************************
.SUBCKT HC00pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHC00     20  30  10  90          INV2
XPK14  2 90  3 90 90 90  0 90 90 90 90 90 90  1 
+     20 90 30 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HCT00pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHCT00    20  30  10  90          INV2T
XPK14  2 90  3 90 90 90  0 90 90 90 90 90 90  1 
+     20 90 30 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HC02pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHC02     20  30  10  90          INV2
XPK14  3  2 90 90 90 90  0 90 90 90 90 90 90  1 
+     30 20 90 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HCT02pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHCT02    20  30  10  90          INV2T
XPK14  3  2 90 90 90 90  0 90 90 90 90 90 90  1 
+     20 90 30 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HC04pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHC04     20  30  10  90          INV1
XPK14  2  3 90 90 90 90  0 90 90 90 90 90 90  1 
+     20 30 90 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HCT04pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHCT04    20  30  10  90          INV1T
XPK14  2  3 90 90 90 90  0 90 90 90 90 90 90  1 
+     20 30 90 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HCU04pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHCU04    20  30  10  90          INV0
XPK14  2  3 90 90 90 90  0 90 90 90 90 90 90  1 
+     20 30 90 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HC05pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHC05     20  30  10  90          INVOD
XPK14  2  3 90 90 90 90  0 90 90 90 90 90 90  1 
+     20 30 90 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HC08pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHC08     20  30  10  90          NINV1
XPK14  2 90  3 90 90 90  0 90 90 90 90 90 90  1 
+     20 90 30 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HCT08pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHCT08    20  30  10  90          NINV1T
XPK14  2 90  3 90 90 90  0 90 90 90 90 90 90  1 
+     20 90 30 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HC14pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHC14     20  30  10  90          INVSMT
XPK14  2  3 90 90 90 90  0 90 90 90 90 90 90  1 
+     20 30 90 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HCT14pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHCT14    20  30  10  90          INVSMTT
XPK14  2  3 90 90 90 90  0 90 90 90 90 90 90  1 
+     20 30 90 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HC32pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHC32     20  30  10  90          NINV1
XPK14  2 90  3 90 90 90  0 90 90 90 90 90 90  1 
+     20 90 30 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HCT32pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHCT32    20  30  10  90          NINV1T
XPK14  2 90  3 90 90 90  0 90 90 90 90 90 90  1 
+     20 90 30 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HC74pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHC74     20  30  10  90          INV1
XPK14 90  2 90 90 90  3  0 90 90 90 90 90 90  1 
+     90 20 90 90 90 30 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HCT74pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHCT74    20  30  10  90          INV1T
XPK14 90  2 90 90 90  3  0 90 90 90 90 90 90  1 
+     90 20 90 90 90 30 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HC86pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHC86     20  30  10  90          NINV1
XPK14  2 90  3 90 90 90  0 90 90 90 90 90 90  1 
+     20 90 30 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HCT86pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHCT86    20  30  10  90          NINV1T
XPK14  2 90  3 90 90 90  0 90 90 90 90 90 90  1 
+     20 90 30 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HC123pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHC123    20  30  10  90          INV1
XPK16  2 90 90 90  3 90 90  0 90 90 90 90 90 90 90  1 
+     20 90 90 90 30 90 90 90 90 90 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HCT123pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHCT123   20  30  10  90          INV1T
XPK16  2 90 90 90  3 90 90  0 90 90 90 90 90 90 90  1 
+     20 90 90 90 30 90 90 90 90 90 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HC132pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHC132    20  30  10  90          INVSMT
XPK14  2 90  3 90 90 90  0 90 90 90 90 90 90  1 
+     20 90 30 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HCT132pck 2 3 1 0
*IN=2, OUT=3, VCC=1, GND=0
XHCT132   20  30  10  90          INVSMTT
XPK14  2 90  3 90 90 90  0 90 90 90 90 90 90  1 
+     20 90 30 90 90 90 90 90 90 90 90 90 90 10 pk14
.ENDS

.SUBCKT HC138pck 2 5 3 1 0
XHC138    20  50  30  10  90      NANDINV
XPK16  2 90 90  5 90 90 90  0 90 90 90 90 90 90  3  1 
+     20 90 90 50 90 90 90 90 90 90 90 90 90 90 30 10 pk16
.ENDS

.SUBCKT HCT138pck 2 5 3 1 0
XHCT138   20  50  30  10  90      NANDINVT
XPK16  2 90 90  5 90 90 90  0 90 90 90 90 90 90  3  1 
+     20 90 90 50 90 90 90 90 90 90 90 90 90 90 30 10 pk16
.ENDS

.SUBCKT HC161pck 2 3 1 0
XHC161    20  30  10  90          INV2
XPK16 90  2 90 90 90 90 90  0 90 90 90 90 90  3 90  1 
+     90 20 90 90 90 90 90 90 90 90 90 90 90 30 90 10 pk16
.ENDS

.SUBCKT HCT161pck 2 3 1 0
XHCT161   20  30  10  90          INV2T
XPK16 90  2 90 90 90 90 90  0 90 90 90 90 90  3 90  1 
+     90 20 90 90 90 90 90 90 90 90 90 90 90 30 90 10 pk16
.ENDS

.SUBCKT HC163pck 2 3 1 0
XHC163    20  30  10  90          INV2
XPK16 90  2 90 90 90 90 90  0 90 90 90 90 90  3 90  1 
+     90 20 90 90 90 90 90 90 90 90 90 90 90 30 90 10 pk16
.ENDS

.SUBCKT HCT163pck 2 3 1 0
XHCT163   20  30  10  90          INV2T
XPK16 90  2 90 90 90 90 90  0 90 90 90 90 90  3 90  1 
+     90 20 90 90 90 90 90 90 90 90 90 90 90 30 90 10 pk16
.ENDS

.SUBCKT HC240pck 2 5 3 1 0
XHC240    20  50  30  10  90      INV3
XPK20  5  2  3 90 90 90 90 90 90  0 90 90 90 90 90 90 90 90 90  1 
+     50 20 30 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 10 pk20
.ENDS

.SUBCKT HCT240pck 2 5 3 1 0
XHCT240   20  50  30  10  90      INV3T
XPK20  5  2  3 90 90 90 90 90 90  0 90 90 90 90 90 90 90 90 90  1 
+     50 20 30 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 10 pk20
.ENDS

.SUBCKT HC244pck 2 5 3 1 0
XHC244    20  50  30  10  90      NINV3
XPK20  5  2  3 90 90 90 90 90 90  0 90 90 90 90 90 90 90 90 90  1 
+     50 20 30 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 10 pk20
.ENDS

.SUBCKT HCT244pck 2 5 3 1 0
XHCT244   20  50  30  10  90      NINV3T
XPK20  5  2  3 90 90 90 90 90 90  0 90 90 90 90 90 90 90 90 90  1 
+     50 20 30 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 10 pk20
.ENDS

.SUBCKT HC245pck 2 5 3 1 0
XHC245   20  50  30  10  90       NINV3
XPK20 90  2 90 90 90 90 90 90 90  0 90 90 90 90 90 90 90  3  5  1 
+     90 20 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 30 50 10 pk20
.ENDS

.SUBCKT HCT245pck 2 5 3 1 0
XHCT245   20  50  30  10  90      NINV3T
XPK20 90  2 90 90 90 90 90 90 90  0 90 90 90 90 90 90 90  3  5  1 
+     90 20 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 30 50 10 pk20
.ENDS

.SUBCKT HC253pck 2 5 3 1 0
XHC253    20  50  30  10  90      NINV3
XPK16  5 90 90 90 90  2  3  0 90 90 90 90 90 90 90  1 
+     50 90 90 90 90 20 30 90 90 90 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HCT253pck 2 5 3 1 0
XHCT253   20  50  30  10  90      NINV3T
XPK16  5 90 90 90 90  2  3  0 90 90 90 90 90 90 90  1 
+     50 90 90 90 90 20 30 90 90 90 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HC273pck 2 3 1 0
XHC273    20  30  10  90          NINV1
XPK20 90  3  2 90 90 90 90 90 90  0 90 90 90 90 90 90 90 90 90  1 
+     90 30 20 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 10 pk20
.ENDS

.SUBCKT HCT273pck 2 3 1 0
XHCT273   20  30  10  90          NINV1T
XPK20 90  3  2 90 90 90 90 90 90  0 90 90 90 90 90 90 90 90 90  1 
+     90 30 20 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 10 pk20
.ENDS

.SUBCKT HC366pck 2 5 3 1 0
XHC366    20  50  30  10  90      INV3
XPK16  5  2  3 90 90 90 90  0 90 90 90 90 90 90 90  1 
+     50 20 30 90 90 90 90 90 90 90 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HCT366pck 2 5 3 1 0
XHCT366   20  50  30  10  90      INV3T
XPK16  5  2  3 90 90 90 90  0 90 90 90 90 90 90 90  1 
+     50 20 30 90 90 90 90 90 90 90 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HC368pck 2 5 3 1 0
XHC368    20  50  30  10  90      INV3
XPK16  5  2  3 90 90 90 90  0 90 90 90 90 90 90 90  1 
+     50 20 30 90 90 90 90 90 90 90 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HCT368pck 2 5 3 1 0
XHCT368   20  50  30  10  90      INV3T
XPK16  5  2  3 90 90 90 90  0 90 90 90 90 90 90 90  1 
+     50 20 30 90 90 90 90 90 90 90 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HC373pck 2 5 3 1 0
XHC373    20  50  30  10  90      NINV3
XPK20  5  3  2 90 90 90 90 90 90  0 90 90 90 90 90 90 90 90 90  1 
+     50 30 20 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 10 pk20
.ENDS

.SUBCKT HCT373pck 2 5 3 1 0
XHCT373   20  50  30  10  90      NINV3T
XPK20  5  3  2 90 90 90 90 90 90  0 90 90 90 90 90 90 90 90 90  1 
+     50 30 20 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 10 pk20
.ENDS

.SUBCKT HC374pck 2 5 3 1 0
XHC374    20  50  30  10  90      NINV3
XPK20  5  3  2 90 90 90 90 90 90  0 90 90 90 90 90 90 90 90 90  1 
+     50 30 20 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 10 pk20
.ENDS

.SUBCKT HCT374pck 2 5 3 1 0
XHCT374   20  50  30  10  90      NINV3T
XPK20  5  3  2 90 90 90 90 90 90  0 90 90 90 90 90 90 90 90 90  1 
+     50 30 20 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 90 10 pk20
.ENDS

.SUBCKT HC595pck 2 5 3 1 0
XHC595    20  50  30  10  90      NINV3
XPK16 90 90 90 90 90 90 90  0 90 90 90 90  5  2  3  1 
+     90 90 90 90 90 90 90 90 90 90 90 90 50 20 30 10 pk16
.ENDS

.SUBCKT HCT595pck 2 5 3 1 0
XHCT595   20  50  30  10  90      NINV3T
XPK16 90 90 90 90 90 90 90  0 90 90 90 90  5  2  3  1 
+     90 90 90 90 90 90 90 90 90 90 90 90 50 20 30 10 pk16
.ENDS

.SUBCKT HC4020pck 2 3 1 0
XHC4020   20  30  10  90          NINV1
XPK16 90 90 90 90 90 90 90  0  3  2 90 90 90 90 90  1 
+     90 90 90 90 90 90 90 90 30 20 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HCT4020pck 2 3 1 0
XHCT4020  20  30  10  90          NINV1T
XPK16 90 90 90 90 90 90 90  0  3  2 90 90 90 90 90  1 
+     90 90 90 90 90 90 90 90 30 20 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HC4040pck 2 3 1 0
XHC4040   20  30  10  90          NINV1
XPK16 90 90 90 90 90 90 90  0  3  2 90 90 90 90 90  1 
+     90 90 90 90 90 90 90 90 30 20 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HCT4040pck 2 3 1 0
XHCT4040  20  30  10  90          NINV1T
XPK16 90 90 90 90 90 90 90  0  3  2 90 90 90 90 90  1 
+     90 90 90 90 90 90 90 90 30 20 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HC4051pck 2 3 4 7 1 0
XHC4051   20  30  40  70  10  90  SWI1
XPK16 90 90  4 90 90  2  7  0 90 90 90 90  3 90 90  1 
+     90 90 40 90 90 20 70 90 90 90 90 90 30 90 90 10 pk16
.ENDS

.SUBCKT HCT4051pck 2 3 4 7 1 0
XHCT4051  20  30  40  70  10  90  SWI1T
XPK16 90 90  4 90 90  2  7  0 90 90 90 90  3 90 90  1 
+     90 90 40 90 90 20 70 90 90 90 90 90 30 90 90 10 pk16
.ENDS

.SUBCKT HC4052pck 2 3 4 7 1 0
XHC4052   20  30  40  70  10  90  SWI1
XPK16 90 90 90 90 90  2  7  0 90 90 90  3  4 90 90  1 
+     90 90 90 90 90 20 70 90 90 90 90 30 40 90 90 10 pk16
.ENDS

.SUBCKT HCT4052pck 2 3 4 7 1 0
XHCT4052  20  30  40  70  10  90  SWI1T
XPK16 90 90 90 90 90  2  7  0 90 90 90  3  4 90 90  1 
+     90 90 90 90 90 20 70 90 90 90 90 30 40 90 90 10 pk16
.ENDS

.SUBCKT HC4053pck 2 3 4 7 1 0
XHC4053   20  30  40  70  10  90  SWI1
XPK16 90 90 90 90 90  2  7  0 90 90 90  3 90  4 90  1 
+     90 90 90 90 90 20 70 90 90 90 90 30 90 40 90 10 pk16
.ENDS

.SUBCKT HCT4053pck 2 3 4 7 1 0
XHCT4053  20  30  40  70  10  90  SWI1T
XPK16 90 90 90 90 90  2  7  0 90 90 90  3 90  4 90  1 
+     90 90 90 90 90 20 70 90 90 90 90 30 90 40 90 10 pk16
.ENDS

.SUBCKT HC4060pck 2 5 3 1 0
XHC4060   20  50  30  10  90      OSC
XPK16 90 90 90 90 90 90  3  0 90 90  2  5 90 90 90  1 
+     90 90 90 90 90 90 30 90 90 90 20 50 90 90 90 10 pk16
.ENDS

.SUBCKT HCT4060pck 2 5 3 1 0
XHCT4060  20  50  30  10  90      OSCT
XPK16 90 90 90 90 90 90  3  0 90 90  2  5 90 90 90  1 
+     90 90 90 90 90 90 30 90 90 90 20 50 90 90 90 10 pk16
.ENDS

.SUBCKT HC4066pck 2 3 4 1 0
XHC4066   20  30  40  10  90      SWI2
XPK14  3  4 90 90 90 90  0 90 90 90 90 90  2  1 
+     30 40 90 90 90 90 90 90 90 90 90 90 20 10 pk14
.ENDS

.SUBCKT HCT4066pck 2 3 4 1 0
XHCT4066  20  30  40  10  90      SWI2T
XPK14  3  4 90 90 90 90  0 90 90 90 90 90  2  1 
+     30 90 90 90 90 90 90 90 90 90 90 90 20 10 pk14
.ENDS

.SUBCKT HC4316pck 2 3 4 7 1 0
XHC4316   20  30  40  70  10  90  SWI3
XPK16  4  3 90 90 90 90 90  0  7 90 90 90 90 90  2  1 
+     40 30 90 90 90 90 90 90 70 90 90 90 90 90 20 10 pk16
.ENDS

.SUBCKT HCT4316pck 2 3 4 7 1 0
XHCT4316  20  30  40  70  10  90  SWI3T
XPK16  4  3 90 90 90 90 90  0  7 90 90 90 90 90  2  1 
+     40 30 90 90 90 90 90 90 70 90 90 90 90 90 20 10 pk16
.ENDS

.SUBCKT HC4538pck 2 3 1 0
XHC4538   20  30  10  90          INVSMT
XPK16 90 90 90  2 90  3 90  0 90 90 90 90 90 90 90  1 
+     90 90 90 20 90 30 90 90 90 90 90 90 90 90 90 10 pk16
.ENDS

.SUBCKT HCT4538pck 2 3 1 0
XHCT4538  20  30  10  90          INVSMTT
XPK16 90 90 90  2 90  3 90  0 90 90 90 90 90 90 90  1 
+     90 90 90 20 90 30 90 90 90 90 90 90 90 90 90 10 pk16
.ENDS
